2 stage OTA. Final aim - use RL agent to design it

* Circuit definition
vin 1 0 dc 0 ac 1
gm1 2 0 1 0 -0.002
r1 2 0 500000.0
c1 2 0 6e-13
cc 2 3 1.25e-11
gm2 3 0 2 0 0.005
r2 3 0 20000.0
c2 3 0 8e-13

.control

***** Analysis command *****
ac dec 10 1e-3 10G

***** Run *****
run

***** Measuring performance metrics *****

* measuring phase margin
let vp_deg = vp(3)*57.29
meas ac phase_margin 
+ FIND vp_deg WHEN vdb(3) = 0

* measuring DC gain
meas ac DC_gain_dB
+ MAX vdb(3) from=1e-3 to=10G 

* measuring UGF
meas ac UGF
+ WHEN vdb(3)=0 CROSS=1

***** Bode plots of vout *****

* Magnitude dB plot for v(3) on log scale
*plot vdb(3) xlog
*+ xlabel 'Frequency in Hz'
*+ ylabel 'Magnitude in dB'
*+ title 'Magnitude plot'

* Phase in degrees plot for v(3) on log scale
*plot {57.29*vp(3)} xlog
*+ xlabel 'Frequency in Hz'
*+ ylabel 'Phase in deg'
*+ title 'Phase plot'

exit ; so that ngspice does not end in interactive mode

.endc
.end
